module a_b(
	input a,
	input b,
	output f
);
	assign f = a ^ b;
endmodule
