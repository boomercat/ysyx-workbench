module alu_ctrl_num(
    input clk,
    input [31:0] instruction,
    output reg [3:0] alu_ctrl
);

// wire [14:0] right_inst;
// assign  right_inst = instruction[14:0];


always @(*) 
begin
  casez (instruction)
    32'b????????????_?????_???_?????_0010111 : alu_ctrl = 4'b0000;     //auipc
    32'b????????????_?????_000_?????_0000011 : alu_ctrl = 4'b0000;     //lb
    32'b0000000?????_?????_000_?????_0110011 : alu_ctrl = 4'b0000;     //add
    32'b????????????_?????_000_?????_0010011 : alu_ctrl = 4'b0000;      //addi: 
    32'b????????????_?????_???_?????_0110111 : alu_ctrl = 4'b0001;    //lui
    32'b????????????_?????_???_?????_1101111 : alu_ctrl = 4'b0000;     //jal   从010->000
    32'b0100000?????_?????_000_?????_0110011 : alu_ctrl = 4'b0010;     //sub
    32'b????????????_?????_000_?????_1100111 : alu_ctrl = 4'b0011;     //jalr
    32'b0000000?????_?????_011_?????_0110011 : alu_ctrl = 4'b0100;      //sltu  和sltiu共用一个
    32'b????????????_?????_01?_?????_0010011 : alu_ctrl = 4'b0100;     ///sltiu -> x[rd] = (x[rs1] < sext(imm))?1:0
    32'b0000000?????_?????_100_?????_0110011 : alu_ctrl = 4'b0101;      //xor ->xori共用
    32'b????????????_?????_100_?????_0010011 : alu_ctrl = 4'b0101;      //xori
    32'b0000000?????_?????_110_?????_0110011 : alu_ctrl = 4'b0110;      //or 跟ori共用
    32'b????????????_?????_110_?????_0010011 : alu_ctrl = 4'b0110;      //ori
    32'b0000000?????_?????_111_?????_0110011 : alu_ctrl = 4'b0111;      //and 跟addi共用一个
    32'b????????????_?????_111_?????_0010011 : alu_ctrl = 4'b0111;      //andi
    32'b0000000?????_?????_001_?????_0110011 : alu_ctrl = 4'b1000;      //sll    跟slli共用一个
    32'b0000000?????_?????_001_?????_0010011 : alu_ctrl = 4'b1000;      //slli
    32'b0000000?????_?????_101_?????_0110011 : alu_ctrl = 4'b1010;      //srl
    32'b0000000?????_?????_101_?????_0010011 : alu_ctrl = 4'b1010;      //srli
    32'b0100000?????_?????_101_?????_0110011 : alu_ctrl = 4'b1010;      //sra    和srai共用一个
    32'b0100000?????_?????_101_?????_0010011 : alu_ctrl = 4'b1001;      //srai
    32'b????????????_?????_010_?????_0010011 : alu_ctrl = 4'b1100;      //slti ->有符号扩展
    32'b0000000?????_?????_010_?????_0110011 : alu_ctrl = 4'b1100;      //slt   有符号扩展
    default: alu_ctrl = 4'b0000;
  endcase
  
end


endmodule